LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY chopper_perder IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=4;
					ADDR_WIDTH	:	INTEGER:=14);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF chopper_perder IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1110","1000","1000","1000","1000","0000","1110","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1000","1101","1101","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","1101","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0111","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0010","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1101","0011","1000","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","1011","0110","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0100","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0011","1000","1110","0011","0011","0011","0011","1010","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","1011","0101","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0011","0011","0011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1011","0001","0001","0001","0001","0001","0001","0001","0001","0101","0100","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","1101","1000","0010","0010","0100","0100","0010","1000","1101","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0111","0100","0100","0111","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1010","0011","0011","0011","0011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","1101","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0011","1101","0001","0001","0001","0001","0001","0001","1011","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0011","0011","0011","0011","0011","0011","0011","1000","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0100","0101","1101","0001","0001","0001","0001","1101","0111","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1100","1101","0001","0001","0001","0001","0001","0001","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0011","0011","0011","0011","0011","0011","1010","0011","0011","0011","1110","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0111","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","1000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","1110","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","1101","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","1110","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1110","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0111","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","1100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","1110","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0011","0011","0011","1000","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0110","1101","1101","0010","0010","0010","0010","0010","1000","1101","1101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0101","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","1110","0000","0000","0000",
     "0000","0000","0000","0000","1101","1101","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0000","0000","0000","0000","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","1101","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","1101","0101","0100","0100","0100","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","1110","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","1000","0000","0000","0000",
     "0000","0000","0000","1101","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1101","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0101","0100","0100","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","1101","0101","0100","0100","0100","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","1110","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","1010","0011","0011","1110","0000","0000",
     "0000","0000","1101","0011","0011","1010","0011","0011","1010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0100","0100","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","1000","0100","0100","0100","0100","0100","0111","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1110","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","1000","0000","0000",
     "0000","0000","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","1000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","0010","0010","0010","0010","1101","0100","0100","0100","0100","0100","0101","0001","0001","0001","0001","0001","0001","0001","0001","1101","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","1101","0000","0000",
     "0000","1000","0011","0011","1101","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","1000","0000","1110","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","1100","1101","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","1101","0110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0010","0010","0010","0010","1101","0101","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","1101","0100","0100","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0011","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","1101","1101","0000",
     "0000","1101","0011","0011","1101","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","1110","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","1101","0001","0001","0001","0001","0101","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","1101","0111","0111","1100","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","0010","0111","0111","1101","0010","0010","0010","0010","1101","0100","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0100","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","1011","0000","0000","0000","1110","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000",
     "0000","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","1000","1110","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","0100","1101","0001","0001","0001","1101","0100","0100","0100","0100","0100","0011","0010","0010","0010","0010","0011","0111","0111","0111","0111","0111","1000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0111","0111","0111","0111","1101","0010","0010","0010","0010","1101","0100","0100","0100","0100","0101","0001","0001","0001","0001","0001","0101","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0000","0000","1110","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1101",
     "0000","0011","0011","0011","0011","0011","0011","0011","1010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1110","1011","0001","0001","0001","0001","0001","0001","0001","0001","1011","0100","0100","0100","0100","1011","0001","0001","0001","0101","0100","0100","0100","0100","0111","0010","0010","0010","0010","0010","1100","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0010","0010","1001","0010","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0100","0100","0100","0100","1101","0001","0001","0001","0001","0010","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1101",
     "0000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0110","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0100","0100","0100","1101","0001","0001","0001","1101","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","0011","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","1001","0100","0111","0111","0111","0111","0111","0101","0111","0111","1101","0010","0010","0010","1010","0101","0100","0100","0100","0111","0001","0001","0001","0001","1011","0111","0100","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0000","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","1000","1000",
     "1110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0010","1011","0001","0001","0001","0001","0101","0100","0100","0100","0100","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","1001","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0011","0010","0010","0010","1101","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0000","1000","0011","0011","0011","0011","0011","0011","1010","0011","0011","0011","0011","1101","0011","0011","0011","1101","1000","1000",
     "0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0100","1000","0010","0010","0010","0011","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0101","0111","0111","0111","0111","0111","0101","0101","0111","0111","0111","0111","1100","0010","0010","0010","1001","0101","0100","0100","0100","0101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1110","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","1101","1000","1000",
     "0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0010","0010","0010","0010","0010","1100","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","1101","1100","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0111","1000","0010","0010","0010","0010","0011","0100","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","1010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","1101","1000","1000",
     "0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0111","0100","0100","0100","0100","1101","0010","0010","0010","0010","1000","1100","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","1000","0100","0100","0100","0100","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1101",
     "0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0100","0100","0100","0100","0100","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0101","0111","1101","0010","0010","0010","0010","0010","0010","0010","0111","0100","0100","0100","0111","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1101",
     "0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0110","0010","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0010","0010","0010","0100","0100","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","1000","1000","1101",
     "0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0110","0100","0100","0100","0100","1101","0010","0010","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","1101","1000","1000","1000",
     "0011","0011","0011","0011","0011","0011","0011","0011","1010","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0100","0100","0100","0100","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","1101","1000","1000","0011",
     "0000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0101","0100","0100","0100","0100","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","0100","0100","0100","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","0000",
     "0000","0011","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","0100","0100","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","1100","0101","0101","0111","0111","0111","0111","0111","0111","0101","0111","0111","0101","0111","0010","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","0100","0100","0100","0100","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1000","0000",
     "0000","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","0100","0101","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0101","0111","0111","0111","0101","0101","0111","0111","0111","0111","0101","0111","0111","0111","0111","0110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0110","0100","0100","0100","0100","0101","0001","0001","0001","1011","0011","0011","1011","0001","0001","0001","0001","0001","0001","0001","1011","1011","1010","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","1101","0011","0011","0011","1101","1000","1000","1000","0000",
     "0000","1010","0011","0011","1101","0011","0011","0011","1101","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0100","0100","0100","0100","0101","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1100","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","0100","0100","0100","0100","0101","0001","0001","0001","0101","0100","0100","0111","0001","0001","0001","0001","0001","0001","0001","1011","1011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","1000","1000","1000","1110","0000",
     "0000","1101","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0010","0101","0011","0001","0001","0001","1011","0100","0100","0100","0100","0101","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","1100","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0010","1001","0010","0010","0010","0010","0010","0010","0010","0010","1010","0100","0100","0100","0100","0101","0001","0001","0001","0111","0100","0100","0100","0001","0001","0001","0001","0001","0001","0001","1011","1101","0011","0011","0011","0011","0011","0011","1010","0011","0011","0011","0011","0011","1010","0011","1000","1000","1000","1000","1000","0000","0000",
     "0000","1000","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0010","0001","0001","0001","0100","0100","0100","0100","0101","1001","0010","0010","0010","0010","0010","0010","0010","0010","1110","1100","0111","0111","0111","0111","0111","0111","0101","0111","0101","0111","0111","0111","0101","0111","0111","0111","0101","0111","0111","0111","0010","1001","0010","0010","0010","0010","0010","0010","0010","1101","0100","0100","0100","0100","0100","0001","0001","0001","0010","0100","0100","0100","0001","0001","0001","0001","0001","0001","0001","1011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","1000","1000","1101","1000","1000","1000","0000","0000",
     "0000","0011","0011","0011","0011","0011","0011","0011","0011","1000","0011","0011","0011","0011","1101","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","0011","0100","0100","0100","0111","0001","0001","0001","0100","0100","0100","0100","0100","1001","0010","0010","0010","0010","0010","0010","0010","1110","1100","0111","0111","0111","0111","0101","0111","0111","0111","0101","0111","0111","0101","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0010","0010","0010","0010","0010","0010","0010","0010","1101","0100","0100","0100","0100","0010","0001","0001","0001","1011","0100","0100","0101","0001","0001","0001","0001","0001","0001","1011","1011","0011","0011","0011","0011","0011","0011","0011","1101","0011","0011","0011","0011","1101","1000","1000","1000","1000","1000","1000","1110","0000","0000",
     "0000","1110","0011","0011","0011","1000","0011","0011","0011","1101","0011","0011","0011","0011","1000","0011","0011","0011","0011","0011","1000","1000","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0001","0001","0001","0111","0100","0100","0100","0100","1000","0010","0010","0010","0010","0010","0010","0011","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0011","0010","0010","0010","0010","0010","0010","1000","0100","0100","0100","0100","1000","0001","0001","0001","0001","0001","1101","0001","0001","0001","0001","0001","0001","0001","1011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1101","1000","1000","1101","1000","1000","1000","0000","0000","0000",
     "0000","0000","1010","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1011","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","1101","0001","0001","0001","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","0010","0010","0101","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0011","1101","0111","0111","0111","0111","0111","0111","0101","0111","0101","0101","0111","0111","1101","0010","0010","0010","0010","0010","0101","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1101","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1000","1000","1000","1000","1101","1000","1000","1000","0000","0000","0000",
     "0000","0000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1101","0001","0001","0001","0001","0001","0001","0001","1101","0100","1101","0001","0001","0001","0001","1000","0100","0100","0100","0100","0010","0010","0010","0010","0010","1001","0101","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","1101","0010","0010","1101","0111","0101","0111","0111","0111","0111","0111","0111","0101","0111","0111","0111","1101","0010","0010","0010","0010","0100","0100","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1101","1000","1000","1000","1000","1000","1000","0000","0000","0000","0000",
     "0000","0000","1110","0011","0011","0011","1101","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0111","0010","0010","0010","0010","0011","0111","0111","0111","0101","0101","0111","0101","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0111","0101","0111","1100","0011","0010","0010","0010","1101","0100","0100","0100","0100","0111","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1101","1000","1000","1101","1000","1000","1101","0000","0000","0000","0000",
     "0000","0000","0000","0011","0011","0011","1000","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0111","0100","0100","0100","0100","1000","0010","0010","0010","1101","0101","0111","0101","0111","0111","0101","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0110","0100","0100","0100","0100","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000",
     "0000","0000","0000","1101","0011","0011","0011","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0100","0100","0100","0100","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0101","0111","1000","0010","0010","0010","0010","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1101","1000","1000","1000","0000","0000","0000","0000","0000",
     "0000","0000","0000","1110","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0100","1000","0010","0010","0010","0010","1101","0111","0111","0111","0111","0111","0111","0111","0010","1000","1101","1000","1000","0011","1101","1101","0010","0010","0010","1101","0111","0111","0111","0111","0111","1101","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1011","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1101","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","1101","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1000","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1100","0100","0100","0100","0100","0110","0010","0010","0010","0010","0010","1101","0111","0101","0111","0111","0101","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","1000","1101","0111","0101","0111","1101","0010","0010","0010","0010","0010","1110","0100","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1011","1011","1011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","0011","0011","1000","1000","1000","1000","1000","1000","1000","1000","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","0010","1101","0111","0110","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","1101","0010","1101","0010","0010","0010","0010","0010","0010","0011","0100","0100","0100","0100","0100","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1011","1011","1011","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1110","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0011","0011","0011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0100","0100","0100","0100","0100","1101","0010","0010","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","1001","0010","0010","0010","1101","0100","0100","0100","0100","0100","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1011","1011","1011","1011","1011","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1110","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0100","0100","0100","0100","0100","0100","1101","0010","0011","1000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","1101","0010","0010","0111","0100","0100","0100","0100","0011","0001","0001","0001","0001","1101","1101","0001","0001","0001","0001","0001","0001","0001","1011","1011","1011","1011","1011","1011","1011","1011","1101","0011","1000","1000","1000","1000","1000","1000","1000","1101","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0011","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0011","0011","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0111","0100","0100","0100","0100","0100","1000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0100","0100","0100","0100","0100","0001","0001","0001","0001","0011","0100","0100","0111","0001","0001","0001","0001","0001","1011","1011","1011","1011","1011","1011","1011","1011","1101","0011","0011","1000","1000","1000","1000","1000","1101","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1000","1000","1000","1000","1000","1000","1000","0011","0011","0011","0011","1101","0001","0001","1011","1000","1101","0001","0001","0001","0001","0001","0001","1101","0100","0100","1101","0001","0001","0001","0001","0001","0001","0101","0100","0100","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0100","0100","1101","0001","0001","0001","1011","0100","0100","0100","0100","1101","0001","0001","0001","0001","1011","1011","1011","1011","1011","1011","1101","1101","0011","0011","1000","1000","1000","1000","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1000","1101","1101","1000","1000","1000","0011","0011","0011","0011","0011","0011","0011","0011","1000","0001","0001","0001","0001","0001","0001","0111","0100","0100","0100","0001","0001","0001","0001","0001","0001","0001","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","1101","0001","0001","0001","0001","1101","0100","0100","0100","0100","1101","0001","0001","0001","1011","1011","1011","0011","0011","0100","0100","0110","1101","0011","0011","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1000","1000","1000","1000","0011","0011","0011","0011","0011","0011","0011","0011","0001","0001","0001","0001","0001","0001","1100","0100","0100","0101","0001","0001","0001","0001","0001","1101","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1001","1101","0001","0001","0001","0101","0100","0100","0100","1101","0001","0001","0001","1011","1011","0011","0011","0100","0100","0100","0100","1101","1000","1000","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0001","0001","0001","0001","0001","0001","0011","0100","0100","1000","0001","0001","0001","1101","1001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0001","1101","0101","1100","1101","0001","0001","0001","1011","1011","1011","0011","1010","0100","0100","0110","0010","1101","1000","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1011","0001","0001","0001","0001","0001","0001","0101","0110","0001","0001","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1000","0001","0001","0001","0001","0001","0001","1011","1011","1011","1101","1000","1000","0011","0011","0010","0011","0011","1000","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1101","1000","1000","1000","1000","1000","1000","1000","1000","1101","1011","0001","0001","0001","0001","0001","0001","0001","0001","1011","1000","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","0001","0001","0001","1011","1011","1011","1011","1101","1000","1000","0011","0011","0011","0011","0011","1000","1000","1000","1000","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0001","0001","1101","1000","1101","1101","1101","0110","0110","0110","0110","1011","0001","0001","0001","0001","0001","0001","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0001","1011","1011","1011","1011","1011","1011","1000","1000","0011","0011","0011","0011","1101","1000","1000","1101","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","1101","1011","0001","0001","0001","1101","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1101","1011","1011","1011","1011","1011","1011","1101","1101","0011","0011","0011","0011","1101","1011","1011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0110","1101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1011","1011","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1110","1000","1101","1010","1010","1010","0011","1101","1101","1110","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1101","1011","1011","1011","1011","1101","0110","0110","1010","1101","1101","1011","1011","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","1010","1010","1010","1010","0110","0110","0110","0110","0110","0110","0110","0110","1011","1011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1110","1101","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1101","1000","1110","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1101","1011","1011","1011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","1000","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1010","1010","1010","1010","1010","1010","0011","0110","0110","0110","0110","1101","1011","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1101","1000","1010","1010","1010","0011","1010","1010","1010","0011","0011","1010","1010","1010","1010","1010","1010","1101","1000","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1101","1011","1000","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1010","1010","1010","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1010","1010","1010","1010","1010","1010","1010","1010","0110","1010","1010","1011","1011","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1101","1010","1000","1010","1010","1010","0011","1010","1010","1010","1010","1010","0011","0011","1010","0011","1010","1010","1101","1010","1010","1000","1101","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1101","1011","0110","0110","0110","0110","0110","0110","0110","0110","0110","1101","1010","1010","1010","1010","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","1010","1010","1010","1010","1010","1010","1010","0011","1010","1101","1011","1011","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1101","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1101","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1101","1011","0110","0110","0110","0110","0110","0110","0110","1101","1010","1010","1010","1010","1010","1010","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1101","0011","0011","1010","1101","1101","0001","0001","0001","1011","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1000","1000","1010","1010","1010","1010","1010","1010","0011","1010","0011","1010","1010","1010","1010","1010","0011","1010","1010","0011","1010","1010","0011","1010","1010","1010","0011","1010","1010","1010","1010","1000","1101","1110","1110","1110","1110","1110","0010","0010","0010","0010","0010","1110","1110","1110","1110","1110","1011","1011","1011","1101","1000","1101","1000","1010","1010","1010","1010","1010","1010","1010","1010","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1011","0010","0010","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1101","1101","0011","0101","1100","0100","0010","1101","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0011","1010","1010","1010","0011","1010","1010","0011","1010","1010","1000","1000","1100","0101","0101","1100","1101","1010","1101","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","0011","1011","1011","1011","1011","1101","1010","1010","1010","0011","1010","1010","1010","1010","1010","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","1110","1110","1110","1110","1101","1010","0011","0101","0101","0101","0101","0101","0101","0101","1100","1101","1010","0011","1010","1010","1010","1010","0011","1010","1010","1010","1010","1010","1010","0011","0011","1010","1010","1101","0101","0101","0101","0101","0101","0101","0101","1100","1101","1010","1101","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1101","1011","1011","1011","1011","1011","1011","1101","1000","1010","1010","0110","1101","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0010","0010","0010","0010","0010","1110","1110","1110","1101","0011","1010","0010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1101","1010","1010","1010","1010","0011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","0010","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1000","1010","1010","0011","1101","1110","1110","1110","1110","1110","1110","1110","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1000","0010","0010","1110","1110","1110","1101","0011","1010","1010","1101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1100","0011","1010","0011","0011","1010","0011","1010","1010","1010","1010","1010","1010","1010","1010","1101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","1010","0011","1010","1010","1011","1101","1110","1110","1110","1110","1101","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","1110","1110","1101","0001","1101","1010","1010","1010","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1101","1010","1010","0011","1010","1010","1010","1010","0011","1010","1010","1010","1010","1010","1100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1010","1010","1010","1010","1011","1011","1011","1101","1101","1101","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","1010","1010","0011","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","1010","0011","1010","0011","1010","1010","1010","1010","0011","1010","1010","1010","1000","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1101","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","1010","1010","1000","0101","0101","0101","0101","0101","0101","0010","0101","0101","0101","0101","0101","0101","0101","1010","1010","1010","0011","1010","1010","1010","1010","1010","0011","1010","1010","1101","0101","0101","0101","0101","0101","0101","1101","1000","0101","0101","0101","0101","0101","1101","1010","0011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","1101","0001","0001","0001","0001","0001","1011","0001","1101","1010","1000","1101","0101","0101","0101","0101","0101","0111","1101","1000","1100","1100","1100","1100","1100","1100","1010","1010","0011","0011","1101","1011","1011","1101","0110","0110","0110","0110","1101","1100","1100","1100","1100","1100","1100","1101","1100","1100","1100","1100","0101","0101","1101","1010","0011","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0001","1101","0011","1010","1000","0101","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","0101","1000","0110","0110","1101","1011","1011","1011","1011","1011","0110","0110","0110","1101","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1010","1010","1010","1010","0001","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","0001","0001","0001","0001","1101","0001","0011","1010","1101","1010","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1101","0110","0110","0110","1011","1011","1011","1011","1011","1011","0110","0110","0110","0110","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","0100","1101","0110","0110","0110","0001","1011","1101","1011","1011","1011","1011","1011","1011","1011","1011","1011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1011","0001","0001","0001","0001","0001","0001","0001","0001","1101","0001","0110","0110","0110","1000","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","0110","0110","0110","0110","1101","1011","1011","1011","1011","1101","0110","0110","0110","0110","0011","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1101","1101","0110","0110","0110","0001","0001","1101","1011","1011","1011","1011","1101","1011","1011","1011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","1011","0001","0001","0001","0001","1011","0001","0110","0110","0110","0110","1101","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1000","1010","0110","0110","0110","0110","1101","1011","1011","1101","0110","0110","0110","0110","0110","0110","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","0010","1000","0110","0110","0110","0110","0001","0001","1011","1011","1011","1011","1011","1101","1011","1011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","1011","1101","0001","0001","0001","0001","0001","0001","0110","0110","0110","0110","1101","0110","1100","1100","1100","1100","1100","1100","1100","1100","1100","0100","0011","0110","0110","0110","0110","0110","0110","0110","1000","0110","0110","0110","0110","0110","0110","0011","1000","1100","1100","1100","1100","1100","1100","1100","1100","0100","1000","0011","0110","0110","0110","0110","0001","0001","1011","0001","1011","1011","1011","1101","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0110","0110","0110","0110","1000","0011","0110","1100","1100","1100","1100","1100","1100","1100","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","1010","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1100","1100","1100","1100","0101","1101","1000","1101","0110","0110","0110","0110","0110","0001","0001","1011","0001","0001","1011","1011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","0001","1010","0110","0110","0110","0110","0110","0110","1101","0010","1100","1100","0101","1101","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0011","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0001","0001","1101","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","1011","1010","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0011","0011","1000","1000","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0001","0001","1101","0001","0001","0001","0001","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","1101","1010","1010","0110","0110","0110","0110","0110","0110","0110","0110","1101","0101","1100","0100","0101","0101","0101","0101","0011","0101","0101","0101","0101","0101","1100","0101","0101","0101","0101","1101","0101","0101","0101","0101","0100","0101","0101","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1011","0001","1101","0001","0001","0001","0001","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","1101","1010","1010","0110","0110","0110","0110","0110","0110","0110","0110","1000","0101","0101","0101","0101","0101","0101","0101","0010","0101","0101","0101","0101","0101","1100","0101","0101","0101","0101","0011","0101","0101","0101","0101","0011","0101","0101","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","1010","1011","0001","1101","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","1101","1000","1010","0110","0110","0110","0110","0110","0110","0110","0110","1101","0101","0101","1100","0101","0101","0101","0101","0010","0101","0101","0101","0101","0101","1100","0101","0101","0101","0101","1100","0101","0101","0101","0101","0011","0101","0101","0100","0110","0110","0110","0110","0110","0110","0110","0110","1010","1010","1011","0001","1011","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","0011","1110","0011","1010","0110","0110","0110","0110","0110","0110","0110","1101","0101","0101","1100","0101","0101","0101","0101","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0101","0010","0110","0110","0011","0110","0110","0110","0110","1010","1010","1101","1101","0001","1011","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","1011","0001","1110","0000","0000","1101","1010","0110","1000","0110","1101","0110","0110","1101","0101","0101","1100","0101","0101","0101","0101","0100","0101","0101","0101","0101","1100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","1100","0101","0101","1101","0110","0110","1101","0110","0110","0110","1101","0011","1000","0000","1101","0001","1011","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","1101","0001","0000","0000","0000","0000","1000","1000","0110","0110","1101","0110","0110","1101","1101","1101","0011","0010","0010","0110","0100","0100","1100","1100","1100","1100","1100","0111","0111","0111","0111","0100","1100","1100","1100","1100","0110","0010","1101","1101","1101","0110","0110","0011","0110","1010","0011","1101","0000","0000","0000","1011","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","1011","0001","0000","0000","0000","0000","0000","0000","0011","1101","1010","0110","0110","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","0110","0110","0110","1101","1000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","1011","0000","0000","0000","0000","0000","0000","0000","0000","1110","0110","0110","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","0110","1010","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0110","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1000","0110","1000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","1011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0110","0011","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","0110","0110","1101","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0110","0110","0110","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1110","1110","1110","1110","1110","1110","1110","1110","1101","1101","1101","1101","1101","1101","1101","1101","0110","0110","1101","1000","0000","0000","0000","0000","0000","0000","0000","1110","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","1011","0001","0011","0000","0000","0000","0000","0000","0000","0000","0000","1010","1101","0110","0110","1101","1101","1101","1101","1101","1101","1101","1101","1110","1110","1110","1110","1110","1110","1110","0011","1110","1110","1110","1110","1101","1101","1101","1101","1101","1101","0110","0110","1010","0011","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","1101","0001","1110","0000","0000","0000","0000","0000","0000","0000","1110","1010","1101","0110","0110","1101","1101","1101","1101","1101","1101","1110","1110","1110","1110","1110","0010","1001","1001","1001","1001","0010","1110","0011","0011","1110","1101","1101","1101","1101","1101","0110","0110","1010","1010","1000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0011","1010","1101","0110","0110","1101","1101","1101","1101","1101","1110","1110","1110","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","1110","1110","1110","1101","1101","1101","1101","0110","0110","1010","0110","1010","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0001","0001","0001","0001","1011","0000","0000","0000","0000","0000","0000","0000","1110","0110","0110","0011","0110","0110","1101","1101","1101","1101","1110","1110","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","1110","1110","1101","1101","1101","0110","0011","1010","0110","0110","0000","0000","0000","0000","0000","0000","0000","1101","0001","1011","0001","0001","0001","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","1000","0110","0110","1010","0110","0110","1101","1101","1101","1110","1110","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1110","1110","1101","1101","1101","0110","1101","0110","0110","0110","1110","0000","0000","0000","0000","0000","0000","0011","0001","1101","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","1011","0001","1000","0000","0000","0000","0000","0000","0000","0000","0011","0110","0110","1101","0110","0110","1101","1101","1101","1110","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1110","1110","1101","1101","0110","1101","0110","0110","0110","0011","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","1110","0000","0000","0000","0000","0000","0000","0000","0110","0110","0110","0101","0011","0110","1101","1101","1110","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","1110","1101","1101","0110","0110","1101","0110","0110","0110","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0001","1101","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","1000","0110","0110","1101","0100","1101","0110","1101","1101","1110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1110","1110","1101","0110","1101","1100","0110","0110","0110","1110","0000","0000","0000","0000","0000","0000","1000","1101","1101","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","0011","0110","0110","0011","1100","1101","0110","1101","0011","0010","1001","1001","1001","1001","1001","1001","1001","1001","0010","1001","1001","1001","1001","0010","1001","1001","1001","1001","1001","1001","0010","1110","0110","0110","1111","0101","1000","0110","0110","0011","0000","0000","0000","0000","0000","0000","0000","0000","1110","1101","1101","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0110","0110","0110","1100","1100","1101","0110","1101","1110","1001","1001","1001","1001","1001","1001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1110","0110","0110","0110","0010","1101","0110","0110","1101","0000","0000","0000","0000","0000","0000","0000","1110","0000","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1011","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","1110","0110","0110","0110","1100","0101","0110","0110","0011","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1110","0110","1101","0110","1101","0101","0110","0110","0011","0000","0000","0000","0000","0000","0000","0000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","1101","0000","0000","0000","0000","0000","0000","0000","1000","0110","0110","1101","0100","1101","0110","0110","0011","0010","1001","1001","1001","1001","0010","1001","1001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","0110","1101","0110","1111","1100","0110","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0001","0001","1000","0000","0000","0000","0000","0000","0000","0000","0110","0110","0110","1101","0100","0011","0110","1101","0110","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1000","0110","1010","1111","0110","0010","1101","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","1101","0000","0000","0000","0000","0000","0000","0000","1110","0110","0110","0110","0010","1100","0110","0110","1101","0110","0010","1001","1001","1001","1001","1001","1001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1101","0110","0110","1111","0110","1101","0011","0110","0110","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0110","0110","0110","1100","1000","0110","0110","1010","0110","1000","1101","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1101","1000","0110","1010","1111","0110","0011","1100","0110","0110","0110","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0110","0110","0110","0110","1100","1101","0110","1111","0110","0110","1000","0101","0010","1101","0010","1001","1001","1001","0010","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1101","0110","0101","0110","1101","1101","0110","0110","0110","1100","0110","0110","0110","0110","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0110","0110","0110","0110","0110","0110","1101","0110","1111","0110","1000","0110","1100","0011","0101","0101","0010","1101","0011","1001","1001","1001","1001","1001","1001","1001","1001","0010","1101","1000","1100","0101","0010","0101","0110","1000","0100","0110","0110","0110","1101","0110","0110","0110","0110","0110","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0110","0110","0110","0110","0110","0110","0110","0011","0110","1111","0110","1101","0110","1101","1100","0101","0101","0101","0101","0111","1100","0100","0110","1000","1101","1000","0100","0101","0101","0101","0101","0101","0101","0010","1101","0110","1100","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0110","0110","0110","0110","0110","0110","0110","1101","0110","0110","0110","1100","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0101","0101","0101","0101","0100","0101","0101","0101","0101","0010","0110","0011","0101","0111","0110","0110","1010","0110","0110","0110","0110","0110","0110","0110","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0110","0110","0110","0110","0110","0110","0110","1101","0110","0110","1101","0101","1101","0110","0011","1100","0101","0101","0111","0101","0101","0101","0101","0010","0101","0101","0101","0101","0101","0101","0101","0101","1100","0011","0110","1000","0101","0101","0110","0110","0011","0110","0110","0110","0110","0110","0110","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","0110","0110","0110","0110","0110","0110","0110","0110","0011","0110","0110","1101","0101","0111","0110","0110","1000","1100","0101","1100","0101","0101","0101","0101","0010","0101","0101","0101","0101","0100","0101","0101","1100","0011","0110","0110","0101","0101","0101","0110","0110","1000","0110","0110","0110","0110","0110","0110","0110","0110","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0110","0110","0110","0110","0110","0110","0110","0110","1010","0110","0110","0100","0101","0101","0010","0110","0110","0011","0100","0111","0101","0101","0101","0101","0010","0101","0101","0101","0101","0100","0101","1101","0110","0110","0110","0010","0101","0101","0101","0110","0110","1000","0110","0110","0110","0110","0110","0110","0110","0110","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0110","0110","0110","0110","0110","0110","0110","0110","0011","0110","0110","0101","0101","0101","0101","1000","0110","0110","0110","1101","0100","0101","0101","0101","0010","0101","0101","0101","0111","1101","0110","0110","0110","0110","0011","1100","0101","0101","0101","0110","0110","0011","0110","0110","0110","0110","0110","0110","0110","1101","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1101","1010","0110","0110","0110","0110","0110","1101","1000","0110","0110","1100","0101","0101","0101","0101","0011","0011","0110","0110","0110","0110","1101","1101","1101","1101","1101","1010","0110","0110","0110","0110","1101","0110","0110","0110","0111","0101","0101","0110","0110","1111","1101","1010","0110","0110","0110","0110","1101","0011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0011","0011","0011","1000","1000","0011","0011","0011","1101","0110","0110","1100","0101","0101","0101","0101","1000","0110","0011","1101","0110","0110","0110","0110","0110","0110","0110","0110","0110","1101","1101","0110","0110","0110","0110","0010","0101","0101","0101","0011","1111","0110","1000","0011","0011","0011","0011","1101","0011","0011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","0011","0011","0011","0011","0011","0011","0011","0011","1000","1111","0110","1100","0101","0101","0101","0101","1000","0110","0110","0110","0110","1101","0010","0011","1000","0010","0010","1100","0101","0101","1101","0110","1111","0110","0110","1000","0101","0101","0101","1000","1111","0110","1101","0011","0011","0011","0011","1101","0011","0011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1000","0011","0011","0011","0011","0011","0011","0011","0110","0110","0110","0101","0101","0101","0101","0101","1000","1111","0110","0110","0110","1000","0111","0101","1100","0101","0101","0101","0101","0101","1101","0110","0110","0110","0110","1000","1100","0101","0101","1101","1111","1101","1000","0011","0011","0011","0011","1101","0011","0011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","0011","0011","1101","1111","1101","1101","0100","1100","0101","0101","0101","1000","0110","0110","0110","0110","1000","0101","0101","0101","0101","0101","0101","0101","0101","0011","0110","0110","0110","0110","0010","1100","0011","1101","1111","1000","1000","1101","1101","0011","0011","1000","1101","0011","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0011","0011","0011","0011","0011","0011","1111","1111","1111","1111","1111","1111","1111","1000","1101","1101","1101","1101","1000","0011","0011","0110","0100","0100","0100","0100","0110","0110","0010","1000","1101","1101","1101","1000","1111","1111","1111","1111","1000","1000","1000","1000","1000","0011","0011","0011","1101","0011","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1101","1000","0011","0011","0011","0011","1101","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1000","1000","1000","0011","0000","1101","0011","0011","1101","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1000","0011","0011","0011","1000","0000","1000","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1000","1000","1110","0000","0000","0000","1101","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1101","1000","1101","0000","0000","1101","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1000","1000","1000","1101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1000","1000","1000","1000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
     "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
	  "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
	  "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
	  "0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000",
	  "0000","0000","0000","0000","0000","0000","0000","0000","0000");
BEGIN 
	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
	   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;