LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Vec_x IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=6;
					ADDR_WIDTH	:	INTEGER:=8);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF Vec_x IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("111111","111110","111101","111100","111011","111010","111001","111000",
												"110111","110110","110101","110100","110011","110010","110001","110000",
												"101111","101110","101101","101100","000001","000010","000011","000100",
												"000101","000110","000111","001000","001001","001010","001011","001100",
												"001101","001110","001111","010000","010001","010010","010011","010100",
												"111111","111110","111101","111100","111011","111010","111001","111000",
												"110111","110110","110101","110100","110011","110010","110001","110000",
												"101111","101110","101101","101100","000001","000010","000011","000100",
												"000101","000110","000111","001000","001001","001010","001011","001100",
												"001101","001110","001111","010000","010001","010010","010011","010100",
												"000010","000011","000100","000101","000110","000111","001000","001001",
												"001010","001011","001100","001101","001110","001111","010000","010001",
												"010010","010011","010100","010101","000000","111111","111110","111101",
												"111100","111011","111010","111001","111000","110111","110110","110101",
												"110100","110011","110010","110001","110000","101111","101110","101101",
												"000010","000011","000100","000101","000110","000111","001000","001001",
												"001010","001011","001100","001101","001110","001111","010000","010001",
												"010010","010011","010100","010101","000000","111111","111110","111101",
												"111100","111011","111010","111001","111000","110111","110110","110101",
												"110100","110011","110010","110001","110000","101111","101110","101101",
												"000010","000011","000100","000101","000110","000111","001000","001001",
												"001010","001011","001100","001101","001110","001111","010000","010001",
												"010010","010011","010100","010101","000000","111111","111110","111101",
												"111100","111011","111010","111001","111000","110111","110110","110101",
												"110100","110011","110010","110001","110000","101111","101110","101101",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000");
BEGIN 
	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
	   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;