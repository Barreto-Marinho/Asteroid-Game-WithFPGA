LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Vec_y IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=6;
					ADDR_WIDTH	:	INTEGER:=8);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF Vec_y IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("010010","010000","001110","001100","001010","001000","000110","000100",
												"000010","000000","111110","111100","111010","111000","110110","110100",
												"110010","110000","101110","101100","010010","010000","001110","001100",
												"001010","001000","000110","000100","000010","000000","111110","111100",
												"111010","111000","110110","110100","110010","110000","101110","101100",
												"101100","101100","101100","101100","101100","101100","101100","101100",
												"101100","101100","101100","101100","101100","101100","101100","101100",
												"101100","101100","101100","101100","101100","101100","101100","101100",
												"101100","101100","101100","101100","101100","101100","101100","101100",
												"101100","101100","101100","101100","101100","101100","101100","101100",
												"010010","010000","001110","001100","001010","001000","000110","000100",
												"000010","000000","111110","111100","111010","111000","110110","110100",
												"110010","110000","101110","101100","010011","010001","001111","001101",
												"001011","001001","000111","000101","000011","000001","111111","111101",
												"111011","111001","110111","110101","110011","110001","101111","101101",
												"010011","010001","001111","001101","001011","001001","000111","000101",
												"000011","000001","111111","111101","111011","111001","110111","110101",
												"110011","110001","101111","101101","010001","001111","001101","001011",
												"001001","000111","000101","000011","000001","111111","111101","111011",
												"111001","110111","110101","110011","110001","101111","101101","101011",
												"010001","001111","001101","001011","001001","000111","000101","000011",
												"000001","111111","111101","111011","111001","110111","110101","110011",
												"110001","101111","101101","101011","010010","010000","001110","001100",
												"001010","001000","000110","000100","000010","000000","111110","111100",
												"111010","111000","110110","110100","110010","110000","101110","101100",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000",
												"000000","000000","000000","000000","000000","000000","000000","000000");
BEGIN 
	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
	   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;