LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Memoria_coseno IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=12;
					ADDR_WIDTH	:	INTEGER:=6);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF Memoria_coseno IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("010000000000","001111111010","001111101010","001111001110",
												"001110100111","001101110111","001100111100","001011111001",
												"001010101101","001001011010","001000000000","000110100000",
												"000100111100","000011010101","000001101011","000000000000",
												"111110010101","111100101011","111011000100","111001100000",
												"111000000000","110110100110","110101010011","110100000111",
												"110011000100","110010001001","110001011001","110000110010",
												"110000010110","110000000110","110000000000","110000000110",
												"110000010110","110000110010","110001011001","110010001001",
												"110011000100","110100000111","110101010011","110110100110",
												"111000000000","111001100000","111011000100","111100101011",
												"111110010101","000000000000","000001101011","000011010101",
												"000100111100","000110100000","001000000000","001001011010",
												"001010101101","001011111001","001100111100","001101110111",
												"001110100111","001111001110","001111101010","001111111010",
												"000000000000","000000000000","000000000000","000000000000");
BEGIN 
	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
	   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;